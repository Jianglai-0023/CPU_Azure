`include "defines.v";
module ALU(

);



endmodule