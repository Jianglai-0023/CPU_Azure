module Decoder(
 input wire         clk,rst,rdy,
 input wire [31:0]  ins,
 input wire         ins_flag,
 input wire [31:0]  pc,
 input wire         pc_bc_flag,
 input wire [31:0]  pc_bc
 //ROB

);








endmodule