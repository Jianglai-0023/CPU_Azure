`include "defines.v";
module ICache(

);

endmodule