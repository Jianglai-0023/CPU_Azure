`include "defines.v";
module LSB(

);

endmodule