`include "defines.v";
module DCache(

);




endmodule